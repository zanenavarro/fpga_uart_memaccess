class uvm_component;
    string name;
    function new(string name);
        this.name = name;
    endfunction
endclass