class uvm_sequencer extends uvm_component;
    function new(string name="uvm_sequencer");
        super.new(name);
    endfunction
endclass