//------------------------------------------------------------------------------
// Module Name    : cmd_execute_tb
// Project        : Latch - UART-Based Register Access System
// Description    : 
//   Structural testbench for verifying the command execution datapath. 
//   Instantiates and ties together the following pipeline of modules:
//
//       uart_rx (stubbed via byte_fifo signals)
//           ↓
//       cmd_parser → cmd_fifo → cmd_dispatcher → register_bank
//
//   Provides a foundation for driver/transaction-based stimulus and response
//   checking. Captures outputs from dispatcher for scoreboard or monitor logic.
//
// Author         : Zane Navarro
// Date Created   : 2025-08-31
// Tool Target    : Vivado / Nexys A7 (Artix-7)
// Synthesizable  : No (Testbench only)
//
// Interfaces     :
//   - Clock/Reset generation (internal in TB)
//   - Byte FIFO interface (stubbed UART RX input)
//   - Command FIFO interface
//   - Dispatcher → Register Bank interface
//   - Dispatcher → TX interface (stubbed for extension)
//
// Revision History:
//   2025-09-08 - Initial version of structural testbench
//------------------------------------------------------------------------------

import cmd_pkg::*;

module cmd_execute_tlb(
    input logic         clk,
    input logic         rst,

    // ---> cmd_parser
    input logic         byte_fifo_valid,
    input logic [7:0]   byte_fifo_data,
    input logic         byte_fifo_rd_en,


    // cmd_dispatcher --->
    output cmd_packet_t cmd_resp_wr_data,
    output logic        cmd_resp_wr_en
);

 

    // cmd parser --> cmd_fifo
    cmd_packet_t cmd_fifo_wr_data;
    logic        cmd_fifo_wr_en;

    // cmd_fifo --> cmd_dispatch
    cmd_packet_t cmd_fifo_rd_data;
    logic        cmd_fifo_rd_en;

    logic        cmd_fifo_valid;
    logic        cmd_fifo_full;
    logic        cmd_fifo_empty;

    // cmd_dispatch <--> register
    logic        reg_read_en;
    logic        reg_write_en;
    logic [7:0]  reg_read_data;
    logic [7:0]  reg_write_data;
    logic [7:0]  reg_addr;


    /////////////////////////////////
    ///////////////////// CMD_PARSER
    cmd_parser cmd_parser (
        .clk(clk),
        .rst(rst),

        // Byte FIFO interface (from uart_rx)
        .byte_fifo_valid(byte_fifo_valid),
        .byte_fifo_data(byte_fifo_data),
        .byte_fifo_rd_en(byte_fifo_rd_en),

        // Command FIFO interface
        .cmd_fifo_wr_en(cmd_fifo_wr_en),
        .cmd_fifo_wr_data(cmd_fifo_wr_data)
        );
    /////////////////////////////////


    /////////////////////////////////
    ///////////////////// CMD_FIFO
    cmd_fifo #(
        .DEPTH(16),
        .ADDR_WIDTH($clog2(16))
    ) cmd_fifo (
        // input
        .clk(clk),
        .rst(rst),

        .wr_en(cmd_fifo_wr_en),
        .wr_data(cmd_fifo_wr_data),

        .rd_en(cmd_fifo_rd_en),

        // output
        .rd_data(cmd_fifo_rd_data),
        .valid(cmd_fifo_valid),
        .full(cmd_fifo_full),
        .empty(cmd_fifo_empty)
    );
    /////////////////////////////////


    /////////////////////////////////
    ///////////////////// CMD_DISPATCH
    cmd_dispatcher cmd_dispatch (
        .clk(clk),
        .rst(rst),

        // input from cmd_fifo
        .cmd_rd_data(cmd_fifo_rd_data),
        .cmd_valid(cmd_fifo_valid),

        //output
        .cmd_rd_en(cmd_fifo_rd_en),
        .mem_addr(reg_addr),

        // output to register file //
        // write
        .mem_write_en(reg_write_en),
        .mem_write_data(reg_write_data),

        // read
        .mem_read_en(reg_read_en),
        .mem_read_data(reg_read_data),
        //////////////////////////////


        // output to RESP FIFO
        .data_out_tx(cmd_resp_wr_data),
        .out_tx_en(cmd_resp_wr_en)
    );

    /////////////////////////////////
    ///////////////////// REGISTER

    register_bank register_bank(
        //input
        .clk(clk),
        .write_en(reg_write_en),
        .read_strobe(reg_read_en),
        .addr(reg_addr),
        .write_data(reg_write_data),

        //output
        .read_data(reg_read_data)
    );
    /////////////////////////////////


endmodule