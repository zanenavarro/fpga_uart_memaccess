class uvm_driver extends uvm_component;
    function new(string name="uvm_driver");
        super.new(name);
    endfunction
endclass