
class mem_access_driver extends uvm_driver;

    virtual mem_access_if vif;
    common_cfg cfg;
    mem_access_transaction cmd_trans;
    mailbox #(mem_access_transaction) seq_mb;


    function new(virtual mem_access_if vif,  common_cfg cfg, mailbox #(mem_access_transaction) seq_mb);
        this.vif = vif;
        this.seq_mb = seq_mb;
        this.cfg = cfg;
    endfunction


    task start();
        int i;
        $display("MEM_ACCESS_DRIVER: Starting mem_access_driver...");

        vif.rx <= 1'b1; // idle state
        @(posedge vif.baud_tick);
    
        for (i = 0; i < cfg.num_sequences; i++) begin
            seq_mb.get(cmd_trans);
            @(posedge vif.baud_tick);
            drive_transaction(cmd_trans);
            @(posedge vif.baud_tick);

        end

    endtask;

    task drive_transaction(mem_access_transaction cmd_trans);
        integer i;
        integer j;
        logic [9:0] data_to_send;

        $display("MEM_ACCESS_DRIVER: Driving cmd_transaction into DUT: cmd_type=%0h, addr=%0h, data=%0h",
            cmd_trans.cmd_type,
            cmd_trans.addr,
            cmd_trans.data);


        // @(posedge vif.baud_tick);
        for (i=0; i<cfg.uart_num_of_byte; i++) begin
        

            // first cmd_type, then cmd_addr, then cmd_data
            data_to_send[8:1] = (i == 0) ? cmd_trans.cmd_type : ((i == 1) ? cmd_trans.addr : cmd_trans.data);
            data_to_send[0] = 1'b0; // start bit
            data_to_send[9] = 1'b1; // stop bit

            $display("MEM_ACCESS_DRIVER: Sending byte %0d: 0x%0h", i, data_to_send[8:1]);

            for (j=0; j<cfg.uart_num_of_bits_tx;j++) begin
                @(posedge vif.baud_tick);
                vif.rx <= data_to_send[j];
            end
            
            @(posedge vif.baud_tick);
        end 
    endtask

endclass