class uvm_monitor extends uvm_component;
    function new(string name="uvm_monitor");
        super.new(name);
    endfunction
endclass