class uvm_scoreboard extends uvm_component;
    function new(string name="uvm_scoreboard");
        super.new(name);
    endfunction
endclass