class reg_access_entry;
    rand logic [7:0] data;

endclass