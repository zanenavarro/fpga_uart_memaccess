class uvm_sequence_itm;
    string name;
    function new(string name="Uvm_sequence_item");
        this.name = name;
    endfunction
endclass